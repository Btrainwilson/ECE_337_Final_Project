// $Id: $
// File name:   tb_FIFO.sv
// Created:     4/19/2018
// Author:      Jackson Barrett
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: test bench for top level block of FIFO design
`timescale 1ns / 10ps

module tb_FIFO();


endmodule

// $Id: $
// File name:   tb_USB_Transmitter.sv
// Created:     4/13/2018
// Author:      Blake Wilson
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: Test Bench USB Timer

module tb_USB_Transmitter();


endmodule

// $Id: $
// File name:   tb_decode.sv
// Created:     2/19/2018
// Author:      Jackson Barrett
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: NRZ decode block test bench
`timescale 1ns / 10ps
module tb_decode ();


endmodule

// $Id: $
// File name:   FIFO.sv
// Created:     4/10/2018
// Author:      Jackson Barrett
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: FIFO buffer for Ethernet-to-USB packet statisitc Collector

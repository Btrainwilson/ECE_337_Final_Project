// $Id: $
// File name:   transceiver_tb_wrapper.sv
// Created:     4/23/2018
// Author:      Luke Upton
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: Testbench wrapper for transceiver

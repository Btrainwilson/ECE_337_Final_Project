// $Id: $
// File name:   tb_rcu.sv
// Created:     2/23/2018
// Author:      Blake Wilson
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: test bench for RCU
`timescale 1ns / 10ps
module tb_rcu ();

	


endmodule

// $Id: $
// File name:   tb_edge_detect.sv
// Created:     2/19/2018
// Author:      Jackson Barrett
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: edge detect test bench for USB reciever
`timescale 1ns / 10ps

module tb_flex_stp_sr ();

endmodule

// $Id: $
// File name:   tb_Byte_Register.sv
// Created:     4/13/2018
// Author:      Blake Wilson
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: test bench for Byte register

module tb_Byte_Register 
();





endmodule

// $Id: $
// File name:   tb_receiver.sv
// Created:     4/17/2018
// Author:      "Stan who drives a Ford"
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: Testbench for receiver side of USB transceiver.


`timescale 1ns / 10ps

module tb_receiver();

	// Define local parameters used by the test bench
	localparam	NORM_CLK_PERIOD		= 10.0 * 100.0 / 96.0; // 10ns * 100 MHz = CLK_PERIOD * 96 MHz.  Everything will be stabilized at 96 MHz after initial syncing)
	localparam	SLOW_CLK_PERIOD		= 10.0 * 100.0 / 96.0 * 1.035;
	localparam 	FAST_CLK_PERIOD		= 10.0 * 100.0 / 96.0 * 0.965;
	localparam 	LINE_CLK_PERIOD		= NORM_CLK_PERIOD;
	localparam DUT_ADDR = 8'b01001100;
    	localparam OTHER_ADDR = 8'b01010010;
    	localparam IN_PID = 8'b01101001;
    	localparam MEH_PID = 8'b00111100;


	// Declare DUT portmap signals
	reg tb_n_rst;
	reg tb_clk;	
	reg tb_d_plus;
	reg tb_d_minus;
	reg tb_is_tx_active;
	reg tb_send_data;
	reg tb_send_nak;
	reg tb_fifo_ready;
	

	// Declare test bench signals
	reg tb_clk_fast;
	reg tb_clk_slow;
	reg tb_line_clk;
	integer tb_test_num;
	integer i;
	integer j;
	
	

	// Clock generation blocks
	always
	begin
		tb_clk = 1'b0;
		#(NORM_CLK_PERIOD/2.0);
		tb_clk = 1'b1;
		#(NORM_CLK_PERIOD/2.0);
	end

	always
	begin
		tb_line_clk = 1'b0;
		#(LINE_CLK_PERIOD/2.0);
		tb_line_clk = 1'b1;
		#(LINE_CLK_PERIOD/2.0);
	end

	// DUT Port map
	receiver DUT(.d_plus(tb_d_plus), .d_minus(tb_d_minus), .clk(tb_clk),
			.n_rst(tb_n_rst), .is_tx_active(tb_is_tx_active),
			.send_data(tb_send_data), .send_nak(tb_send_nak),
			.fifo_ready(tb_fifo_ready));

	// Test vector struct
	//typedef struct
	//{
	//	reg first_bit; // Bit prior to encoded message
	//	reg [7:0] unencoded;
	//} testVector;


	task resetDUT;
	begin
		// Power-on reset of DUT
		tb_n_rst = 1'b0;
		@(negedge tb_clk);
		@(negedge tb_clk);
		tb_n_rst = 1'b1;
		@(negedge tb_clk);
		@(negedge tb_clk);

	end
	endtask

	task send_byte;
		input [7:0] line_byte;
	begin
		for(i = 0; i < 8; i += 1)
		begin
			send_bit(line_byte[i]);
		end

	end
	endtask

	task send_bit; // Sends encoded bit using specified clocking rate.
		input bit_in;
	begin
		if(bit_in == 1'b0)
		begin
			tb_d_plus = ~tb_d_plus;
			tb_d_minus = ~tb_d_plus;
			for(j = 0; j < 8; j++)
			begin
				@(negedge tb_line_clk);
			end
		end
		else
		begin
			tb_d_plus = tb_d_plus;
			tb_d_minus = ~tb_d_plus;
			for(j = 0; j < 8; j++)
			begin
				@(negedge tb_line_clk);
			end
		end
	end
	endtask

	task send_eop;
	begin
		tb_d_plus = 0;
		tb_d_minus = 0;
		for(j = 0; j < 16; j++)
		begin
			@(negedge tb_line_clk);
		end
		tb_d_plus = 1;
		tb_d_minus = 0;
		for(j = 0; j < 8; j++)
		begin
			@(negedge tb_line_clk);
		end
		
	end
	endtask

	initial  // HEY!!! THE TEST'S DOWN HERE
	begin
	// initialize yo crap
	tb_d_plus = 1;  // Idle
	tb_d_minus = 0;
	tb_is_tx_active = 0;
	tb_fifo_ready = 0;

	// power-on reset
	resetDUT();
	
	// Test 1: Send sync byte, correct PID,DUT_address.  Will send nak (fifo not ready).
	tb_test_num = 1;
	send_byte(8'b10000000);
	send_byte(IN_PID);
	send_byte(DUT_ADDR);
	// Should wait until eop is processed now.
	@(negedge tb_clk);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 0;
	tb_d_minus = 0;
	// send_nak should pulse
	@(posedge tb_send_nak);
	assert(tb_send_nak == 1)
            $info("Test %d: PASS - Send nak properly triggered", tb_test_num);
        else
            $error("Test %d: FAIL - Send nak did not properly trigger", tb_test_num);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 1;
	tb_d_minus = 0;
	// send_nak should deassert
	assert(tb_send_nak == 0)
	    begin
            $info("Test %d: PASS - Send nak properly deasserted", tb_test_num);
	    $info("Test %d: Accepts correct PID, Address, and broadcasts nak (fifo not ready)", tb_test_num);
	    end
        else
            $error("Test %d: FAIL - Send nak did not properly deassert", tb_test_num);

	// Test 2: Send sync byte, correct PID,DUT_address.  Will send data (FIFO's BODY IS READY).

//&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&%%%&&&&&%%%%&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&%%%%%&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&%%%%%%&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&@@&&&&&&&&&&&&&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&@@@@&&&&&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&
//&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&%%%&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&%%%%%%%%&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&%%%%%%%%%%%%%%%%&&&&&&&&&&&&%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&%%%%%%%%%%%%%%%%%&&&&&&&&&&%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&%%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&%%%%%%&&%%%%%&&&&&%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&%%%%%%%%%%%&&&&&&&%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&%%%%%%%%&&&&&&&&&%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&%%&&&&&&&&&&&%%%%%%&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&%%%%%&&&&&&&&&&&&%%%%&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&%%%%%%%%&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@@@@@@@@@@@@&&&%%%%%%%%%%%%&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%%%%%%%%%&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&@@@@@@@@@@@@@@@&&&&%%%#((//////////((((((((######%%%%%%%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&%%%%%%%&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@@@@@@@@@@&&&%#(((////*******************////////((((###%%%%&&&&&&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&%&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@@@@@@@@@&%###(/////************************/////////(((####%%%%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@@@@@&&%##(////*****************************////////////((((((((((####%%&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@@@@%##((//////********************************/////////(((((((((((((((##%%%&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@@@&%##(//////*********************************/////////((((((((((((((#####%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&@@@@@@@@@@%#(((/////**********************************/////////(((((((((((((######%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@@@&%#((//////**********************************///////////(((((((((((####%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@&%(((//////**********************************///////////(((((((((((####%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@&(((//////*******************************///////////////((((((((######%%%%&&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@&%#(////////********************************///////////////(((((((######%%%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@@@@@@@&%#(////////**********************************/////////////(((((((######%%%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@(////////**********************************////////////((((((((######%%%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&&&&&&&&&%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&%&&@@@@@@@@%#(////////**********************************////////////((((((((########%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&%&&@@@@@@@@%#(//////************************************/////////////(((((((((######%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&&&&&&%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&@@@@@@@@%((/////***************************************////////////((((((((#######%%%&&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%&&&&%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&%&%%%%&&&@@@@@@@&%(/////***************************************//////////////(((((((#######%%%%%&&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&%%%%&&&&&@@@@@&%(////************************************////////////////////((((((#########%%%%&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&&&%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&@@@@(///*******************************////////////////((((((#((((((((((############%%%&@@@@@@@@@@@@@@@@@@@@@@@@@@@@@@&&&&%%&&&%%&&%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&@@@/////*******////************////*/////////((((((((((#######################%#####%%%&&@@@@@@@@@@@@@@@@@@@@@@&&&&&@@&&&%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&%%&&&&@&&%(((((///////////////////////////////(((((####%%%&&&&&&&&%%%%%%%%%%%%#####%###########%%&&&&@@@@@@@@@@@@@@@@&&%%%%%%%&&&%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&%%&&&&&&&%##%%%%##########((((((((//////////(((####%%%%&&&&&&&&&&&%%%%%%%%%%%%%%%%%%%%%##########%%%%&@@@@@@@@@@@@@@@&&%%%%&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&@&&%#%%%%%%&&&&&%%%%####(((((////////(((####%%%&&&&&&&&&&&&&&&%%%%%%%%%%%%%%%%%%%###########%%%&&@@@@@@@@@@@@&&&%%%%%&%%##%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&%&&&@@@@&%%%%%%&&&&&&&&@@&&&&%%%##(((((((((###%%%%&&&&&@&&&%%%%%%&@@@@@&&&&&%%%%%%%%%%#############%%&&@@@@@@@@@@@&&&%%%%%&&%###%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&@@@&%%%%%&&&&%%%&&&&@@@@&&&%#(////////((###%&&&&&&%%((//#&&&@@@&%%#%&&&&%%%####################%%&&&@@@@@@&&&&&&%%%%%%&%##(#%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&@&&%%%%&&&&###&&&&@@@&&&&(//***///((#%%%&&&&&&%#//**(%&&@@@&%%##%%%%%%####(((((############%%&@@@@@@@&&&&&&&%%%%%%&%##(#%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&##%%%&%(///(%&@@@@&%%%%%#(//**////((###%%%####((/////(######((########(((((((((((((((#######%&&&@@@&&&&&&%%%%%%###%%##(#%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&%%#((####(((///(#######(((((///*////((((#####((((((((((((((((######(((((//////((((((((((#######%%%%&&&&&%%&&&&&&&%%%###(((#%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&%%((((((((((((((((((((###((/////////(((((((#(((((((((((##########(((/////////(((((((((((#######%%%%%%%%%%%&&&&&&&%%%###(((#%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%##(//////((((((((###(((((/////////(((((((((((((((((///(((((((((/////****/////(((((((((((########%%%%%%%%%%%&&&&&&&%%###(((%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((//////////(((((((//////(////////((((((((((((////////////////////******//////(((((((((###%%%##%%%%%%%%%%#%%&&&&&%##(((((#%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((///////////////////////////////((((((((((//////////////////***********//////(((((((((###%%%%%%%%%%%%%%%##%&&&&&%(((((((#%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#/////******//////////////////////(((((((((((///////////////*************///////((((((#####%%%%%%%%%%%%%%##%&&&&&%((((((((%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%(/////*******//////////////////////((((((((((((((//////*/////***********///////(((((((#####%%%%%%%%%%%%%%%%%&%%###((((((##%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#(/////**************///////***/////(((((###((((((((/*****************////////((((((((#####%%%%%%%%%%%%%%%%%%%((//(#((//(%%&%%&%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#(////////*********////////**,***///(((((((((((((((((//*************//////////(((((((#####%%%%%%%%%%%%%%%%%%#(((//((((/(%%%%%&%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#(////////*********////////******/////(((((((/(((((#(////**********///////////((((((######%%%%%%%%%%%%%%%%%%#(((//(((((#%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#(////////********/////////////////(((((((////(((((##((///*******//////////(((((((#######%%%%%%%%%%%%%%%%%%%#(((///(((#%%&&&%%&&&&%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#(////////////***/////((((((///((((###############%%%##(/////**/////////((((((((#######%%%%%%%%%%%%%%%%%%%%##(((//((##%%&&&%%%%&&&%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#(///////////////////(#####((((((##%%%%%&&&&&%%%%%%&&%%(////////////////((((((((#######%%%%%%%%%%%%%%%%%%%%##((((((#%%%&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#(((/////////////////(#%&&&&%%%%%%%&&&&&&&&&&&&&&&&%%##(((///////////((((((((((########%%%%%%%%%%%%%%%%%%%%%##%%%%%%%%%&%%%%&%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((////////((((((((((((######%%%&&&&&&&%%%%########((((((((((//((((((((((((##########%%%%%%%%%%%%%%%%%%%%%%%&&&&&%&&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((//((((((((((((((((((((((((###%%%%%%%###########(((((((((((((((((((((((((##########%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((((((//((##(((((((((((((((((((((((((((((((((((((#######((((((((((((((((((###########%%%%%%%%%%%%%%%%%%%%%%%&&&&&%%%&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%##((((((((#(((((((((///////////////////((((((((((((((######(((((((((((((((((#########%%%%%%%%%%%%%%%%%%%%%%%&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%##((((((((((((((((((///((///////////(((((((((((((((((####(((((((((((((((((((#########%%%%%%%%%%%%%%%%%%%%%%%&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%###(((///(((((((((((((((((((((((((((####%%%%%%%%%%%%%%%%###(((((((((//((((((###(((#####%%%%%%%%%%%%%%%%%%%%%%%&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((///////(((((((#%%%%%%%%%%%%%%%%%&&&&&%%%%&&&&&&&&&&%##((((((((////(((((##(((((####%%%%%%%%%%%%%%%%%%%%%&&&&%%&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((/////////((((((#%%%%%#######%%%%%##########%%%%%%%%#((((((((((////(((((##(((((####%%%%%%%%%%%%%%%%%%%%%&&&&%%&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((//////////////(((((((((((/////////(((((((((#####(((////(////////(((((((((((((##%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&%%%%&&%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((///////////////(((((((////*****//((((((((((####((/////////////((((((((((((((##%%%%%%%%%%%%%%%%%%%%%%##%%%&&&&&&%%%%&&%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#(((//////////////(((((((((/////((((#########((((//////////////((((((#((((((###%%%%%%%%%%%%%%%%%%%%%%###%%&@@@@@@&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((((/////////////((((((((((((((###(((((((((((((///(////////((((((((((((((###%%%%%%%%&&&&%%%%%%%%########%&@@@@@@&&&&&%%%%%%%%%%%%%%%%%%%%%%%&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((((/////////////(((((((((((((((((((((/(((((////(((((////(((((((((((((((##%%%%%%%%%%&&&&%%%%%%%%########%&@@@@@@@&&&&%%%%%%%&&&%%%%%%%%%%%%&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%##(((//////////////////////(((((/////////////((((((((///((((((((((((#####%%%%%%%%%&&&&&&%%%%%%#####(####%&@@@@@&&&&&&&&%%%%%&&&&&%%%%%%&&&&%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%##((//////////////////////////////////////(((((((///(((((((((((######%%%%%%%%%%%&&&&&&%%%#####(((#####%&&&&&&&&&&&&&&&&&%%&&&&&%%%%%%&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%#((((/////////////////////////////////////(((((((((((((((((########%%%%%%%%%%%&&&&&&&%%%#####(((###%%&&&&&&&&&&&&&&&&&&&%%&&&&&%%%%&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%##((((//////////////////////////////////////((((((((((((#######%%%%%%&&&&&&&&&&&&&&%%############%%%&&&&&&&&&&&&&&&&&&&&%%%&&&%%%&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%##(((((////////////*******////////////////(((((((##########%%%%%&&&&&&&&&&&&&&%%%%############%&&&&&&&&&&&&&&&&&&&&&&&&%%&&&%%%%%&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%###((((//////////**********///////////////(((((#########%%%%%%&&&&&&&&&&&&&&&&%%%#############%&&&&&&%%%%%%%%&&&&&&&&&&&&%%%%%%%%%&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%##(((////////////////***//////////(((((((#####%%%%%%%%%%&&&&&&&&&&&&&&&&&%%###############%&&%%%%%%%%%%%%%%%%%&&&&&&&&%%%%%%%%%%%&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&%%%##((/////((((((((((///(/////(((((((((###%%%%%%%%%%&&&&&&&&&&&&&&&&&&%%%%###############%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&%%&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&%%%###((////((((((((((((((((///((((((((###%%%%&&&&&&&&&&&&&&&&&&&&&&&&%%%%##############%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&%%&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&%%%#((((((((((((((((((((((((((((####%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&%%##############(##%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&%%%&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&%%##((((((((########((((((####%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&%%%%#########(((((((#%%%%%%%%%%%%%##%%%%%%%%%%%%%%&&&&%&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&%%%###(((#######((########%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&%%%%########((((((((##%%%%%%%%%%%%%###%%%%%%%%%%%%%&&&%%%&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&%%%%%######(#####%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&%%%########(((/////(###%%%%%%%%%%%%%%%%##%%%%%%%%%%&&&%%%%%%%%%%&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&%%%%%%######%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&%%%########(((//////(##%%%%%%%%%%%%%%%####%%%%%%#%%%&&&&&&&&&&&&%%%%%&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&%%%%%%%%%%%%%%%%%%&&&&%%%%%%%%&&&&&&&&&&&&&&&&&%%%%#####(((////*****/(#%%%%%%%%%%%%%######%%%###%%%%%&&%%%%%&&&&&&&&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&%%%%%%%%&&&&&&&&&%%%%%%%%%%%%&&&&&&&&&&&&&&&&%%%%%%###((((//********/(#%%%%%%%%%%%%%%####%%%%###%%%%&&&%%%%%%%%%%%%%&&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&%%%%%%#####(((//******,**/##%%%##%######%%####%%%%#%%%%%%&&%%%%%%%%%%%%%%%&&&&&
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&&&&&&&&%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&%%%%%%%####((////****,,,*//#%%%%%%%%%%%%%%%%%%%%%%%%%##%%&&%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&%%%&%%%#%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&%%%%%%%%#####((//****,,,,,*(###%%%%%%%####%%%%%%%%%%%%##%%%%&%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&&&&&&&%%&&&%##%%%%%%%%%%%%%%%%&&&&&&&&&&&&%%%%%%%%####(((///***,,,,,,/#%%%%%#%%%%####%%%%%%%%%%%%##%%%&&%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&%&&&&&&&&%%%%(/((###%%%%%%%%%%%%&&&&&&&&&%%%#########((((//****,,,,,*/####%%%%%%%%%%%%#%######%%%%%#%%&&%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&%%%%%%%%%%%%&&&&&&&&&&&&&&&&&&&%%%%%%%%%#***(#######%%%%%%%&&&%%%##########((((((////***,,,,,**/##############%%###############%%&&%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&%%%%%%%%%%#*,,*(#######%%%%%%%%%######(((((((((((/////***,,,,,,**(##############################%%%&%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&%%%%%%%%%%%%#*,,,,*(########%##((///((((/((/////////*****,,,,,,,*((##########%%%#%%%%%%######%####%&&&%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&%/,,,,,,**(#####(/*******/////////********,,,,,,,,,*(################################%%&&%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&%%%%%%%%%%%%%%%%%%&&&%(,,,,,,**/(((//*,,,,********************,,,,,,,,,*/#################################%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&&%%%%%%%%%%%%%%%%%&&&&&**,,,,*****,,,,,,,,,,,,,,,,*****,,,,,,,,,,,,,,**/#############################%###%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&%%%%%%%%%%%%%%%%%%%%&&&&&&//,,,******,,,.,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,//(#################################%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&%#//*/(#((//*,.........,,,,,,,,,,,,,,,,,,,,,,,,/((##################################%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&%%(//(##/////(/,,........,,,,,,,,,,,,,,,,,,,,,,*(##%#%%%###########################%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&%#(((#%%#((/(#(**.........,,,,,,,,,,,,,,,,,,,,,/#%%%%#################%%%%%%####%%#%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%
//%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%&&&%%%%%%%%%%%%%%%%%%%%%%%%&&&&&&&&&&%%%####%&%###((((//*,.......,,,,,,,,,,,,,,,,,,,*/###################%%%%%%%%%########%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%%


	resetDUT();
	tb_fifo_ready = 1;
	tb_test_num += 1;
	send_byte(8'b10000000);
	send_byte(IN_PID);
	send_byte(DUT_ADDR);
	// Should wait until eop is processed now.
	@(negedge tb_clk);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 0;
	tb_d_minus = 0;
	// send_data should pulse
	@(posedge tb_send_data);
	assert(tb_send_data == 1)
            $info("Test %d: PASS - Send data properly triggered", tb_test_num);
        else
            $error("Test %d: FAIL - Send data did not properly trigger", tb_test_num);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 1;
	tb_d_minus = 0;
	// send_data should deassert
	assert(tb_send_data == 0)
	begin
            $info("Test %d: PASS - Send data properly deasserted", tb_test_num);
	    $info("Test %d: Accepts correct PID, Address, and broadcasts data (fifo is ready)", tb_test_num);
	end
        else
            $error("Test %d: FAIL - Send data did not properly deassert", tb_test_num);

	// Test 3: Send sync byte, incorrect PID,DUT_address.  Will send nak (fifo ready, but PID incorrect).
	resetDUT();
	tb_fifo_ready = 1;
	tb_test_num += 1;
	send_byte(8'b10000000);
	send_byte(MEH_PID);
	send_byte(DUT_ADDR);
	// Should wait until eop is processed now.
	@(negedge tb_clk);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 0;
	tb_d_minus = 0;
	// send_nak should pulse
	@(posedge tb_send_nak);
	assert(tb_send_nak == 1)
            $info("Test %d: PASS - Send nak properly triggered", tb_test_num);
        else
            $error("Test %d: FAIL - Send nak did not properly trigger", tb_test_num);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 1;
	tb_d_minus = 0;
	// send_nak should deassert
	assert(tb_send_nak == 0)
	begin
            $info("Test %d: PASS - Send nak properly deasserted", tb_test_num);
	    $info("Test %d: Accepts incorrect PID, correct Address, and broadcasts nak (fifo is ready)", tb_test_num);
	end
        else
            $error("Test %d: FAIL - Send nak did not properly deassert", tb_test_num);

	// Test 4: Send sync byte, correct PID,incorrect address.  Will send nothing (fifo ready, but command not addressed to device).
	resetDUT();
	tb_fifo_ready = 1;
	tb_test_num += 1;
	send_byte(8'b10000000);
	send_byte(IN_PID);
	send_byte(OTHER_ADDR);
	// Should wait until eop is processed now.
	@(negedge tb_clk);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 0;
	tb_d_minus = 0;
	// send_data and send_nak shouldn't pulse (check for a couple clock cycles after broadcasting eop)
	@(negedge tb_clk);
	assert(tb_send_nak == 0 && tb_send_data == 0)
            $info("Test %d: PASS - nak and/or data lines did not trigger - window 1", tb_test_num);
        else
            $error("Test %d: FAIL - nak and/or data lines did trigger - window 1", tb_test_num);
	@(negedge tb_clk);
	assert(tb_send_nak == 0 && tb_send_data == 0)
            $info("Test %d: PASS - nak and/or data lines did not trigger - window 2", tb_test_num);
        else
            $error("Test %d: FAIL - nak and/or data lines did trigger - window 2", tb_test_num);
	@(negedge tb_clk);
	assert(tb_send_nak == 0 && tb_send_data == 0)
            $info("Test %d: PASS - nak and/or data lines did not trigger - window 3", tb_test_num);
        else
            $error("Test %d: FAIL - nak and/or data lines did trigger - window 3", tb_test_num);
	tb_d_plus = 1;
	tb_d_minus = 0;
	// send_nak should deassert
	@(negedge tb_clk);
	assert(tb_send_nak == 0 && tb_send_data == 0)
            $info("Test %d: PASS - nak and/or data lines did not trigger - window 4", tb_test_num);
        else
            $error("Test %d: FAIL - nak and/or data lines did trigger - window 4", tb_test_num);
	@(negedge tb_clk);
	assert(tb_send_nak == 0 && tb_send_data == 0)
            $info("Test %d: PASS - nak and/or data lines did not trigger - window 5", tb_test_num);
        else
            $error("Test %d: FAIL - nak and/or data lines did trigger - window 5", tb_test_num);

	// Test 5: Send sync byte, correct PID,correct address (without resetting DUT).  Will send data (fifo ready, but command not addressed to device).
	tb_fifo_ready = 1;
	tb_test_num += 1;
	send_eop;
	send_byte(8'b10000000);
	send_byte(IN_PID);
	send_byte(DUT_ADDR);
	// Should wait until eop is processed now.
	@(negedge tb_clk);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 0;
	tb_d_minus = 0;
	// send_data should pulse
	@(posedge tb_send_data);
	assert(tb_send_data == 1)
            $info("Test %d: PASS - Send data properly triggered", tb_test_num);
        else
            $error("Test %d: FAIL - Send data did not properly trigger", tb_test_num);
	@(negedge tb_clk);
	@(negedge tb_clk);
	tb_d_plus = 1;
	tb_d_minus = 0;
	// send_data should deassert
	assert(tb_send_data == 0)
	begin
            $info("Test %d: PASS - Send data properly deasserted", tb_test_num);
	    $info("Test %d: Accepts correct PID, Address, and broadcasts data (fifo is ready)", tb_test_num);
	end
        else
            $error("Test %d: FAIL - Send data did not properly deassert", tb_test_num);
	
	end
endmodule

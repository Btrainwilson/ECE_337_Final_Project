// $Id: $
// File name:   tb_shift_register.sv
// Created:     2/23/2018
// Author:      Blake Wilson
// Lab Section: 337-02
// Version:     1.0  Initial Design Entry
// Description: shift register test bench
